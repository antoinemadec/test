/******************************************************************************
  FILE : reset_if.sv
 ******************************************************************************/
interface reset_if (input clock, output logic resetN);
endinterface : reset_if
