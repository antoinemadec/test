library IEEE ;
use IEEE.STD_LOGIC_1164.all ;

package	constants is
        type TPicoType is ( pbtI, pbtII, pbt3, pbtS ) ;
	constant PicoType  : TPicoType := pbt3 ;
	CONSTANT ADDRSIZE  : natural := 10;
	CONSTANT INSTSIZE  : natural := 18;
	CONSTANT JADDRSIZE : natural := 11;
	CONSTANT JDATASIZE : natural := 9;
end package ;


library IEEE ;
use IEEE.STD_LOGIC_1164.all ;
use IEEE.STD_LOGIC_ARITH.all ;
use IEEE.STD_LOGIC_UNSIGNED.all ;

library unisim ;
use unisim.vcomponents.all ;

use work.constants.all;

entity prog_ram is
    port ( 
        clk         : in  std_logic ;
        address     : in  std_logic_vector( ADDRSIZE - 1 downto 0 );
        instruction : out std_logic_vector( INSTSIZE - 1 downto 0 );
        ext_addr    : in  std_logic_vector( JADDRSIZE - 1 downto 0 );
        ext_data    : in  std_logic_vector( JDATASIZE - 1 downto 0 );
        ext_write   : in  std_logic ;
        out_data    : out std_logic_vector( JDATASIZE - 1 downto 0 )
    ) ;
end entity prog_ram ;

architecture mix of prog_ram is

    attribute INIT_00 : string ;
    attribute INIT_01 : string ;
    attribute INIT_02 : string ;
    attribute INIT_03 : string ;
    attribute INIT_04 : string ;
    attribute INIT_05 : string ;
    attribute INIT_06 : string ;
    attribute INIT_07 : string ;
    attribute INIT_08 : string ;
    attribute INIT_09 : string ;
    attribute INIT_0A : string ;
    attribute INIT_0B : string ;
    attribute INIT_0C : string ;
    attribute INIT_0D : string ;
    attribute INIT_0E : string ;
    attribute INIT_0F : string ;
    attribute INIT_10 : string ;
    attribute INIT_11 : string ;
    attribute INIT_12 : string ;
    attribute INIT_13 : string ;
    attribute INIT_14 : string ;
    attribute INIT_15 : string ;
    attribute INIT_16 : string ;
    attribute INIT_17 : string ;
    attribute INIT_18 : string ;
    attribute INIT_19 : string ;
    attribute INIT_1A : string ;
    attribute INIT_1B : string ;
    attribute INIT_1C : string ;
    attribute INIT_1D : string ;
    attribute INIT_1E : string ;
    attribute INIT_1F : string ;
    attribute INIT_20 : string ;
    attribute INIT_21 : string ;
    attribute INIT_22 : string ;
    attribute INIT_23 : string ;
    attribute INIT_24 : string ;
    attribute INIT_25 : string ;
    attribute INIT_26 : string ;
    attribute INIT_27 : string ;
    attribute INIT_28 : string ;
    attribute INIT_29 : string ;
    attribute INIT_2A : string ;
    attribute INIT_2B : string ;
    attribute INIT_2C : string ;
    attribute INIT_2D : string ;
    attribute INIT_2E : string ;
    attribute INIT_2F : string ;
    attribute INIT_30 : string ;
    attribute INIT_31 : string ;
    attribute INIT_32 : string ;
    attribute INIT_33 : string ;
    attribute INIT_34 : string ;
    attribute INIT_35 : string ;
    attribute INIT_36 : string ;
    attribute INIT_37 : string ;
    attribute INIT_38 : string ;
    attribute INIT_39 : string ;
    attribute INIT_3A : string ;
    attribute INIT_3B : string ;
    attribute INIT_3C : string ;
    attribute INIT_3D : string ;
    attribute INIT_3E : string ;
    attribute INIT_3F : string ;
    attribute INITP_00 : string ;
    attribute INITP_01 : string ;
    attribute INITP_02 : string ;
    attribute INITP_03 : string ;
    attribute INITP_04 : string ;
    attribute INITP_05 : string ;
    attribute INITP_06 : string ;
    attribute INITP_07 : string ;
begin
	I18: IF PicoType = pbt3 GENERATE
  	  attribute INIT_00 of bram : label is "000054024044501340545033405250464050505D404C5084404D0072008B0001" ;
	    attribute INIT_01 of bram : label is "A1008001002F002F002F002FC2BAC0B99210028001000000006A40020080008B" ;
	    attribute INIT_02 of bram : label is "0FFF40025C23E100C001002F002F002F002FC2BAC0B99210028001FF00FE5C16" ;
	    attribute INIT_03 of bram : label is "4110C010007292004010C01000724213C2134210C01000720078A0005C30CF01" ;
	    attribute INIT_04 of bram : label is "91004010C01000724113C1134110C010007200784002C27F006AC17E4113C113" ;
	    attribute INIT_05 of bram : label is "C010007200784002D210006A92004010C01000724213C2134210C01000720078" ;
	    attribute INIT_06 of bram : label is "400AC0034003506A200140024002C100006A91004010C01000724113C1134110" ;
	    attribute INIT_07 of bram : label is "4078B0004F20CF034F0350782F014F02A000C0034003507220014002406AB000" ;
	    attribute INIT_08 of bram : label is "8E00CE08CF090E800F0643E9C008C0090000008B0002006AA000548020024002" ;
	    attribute INIT_09 of bram : label is "B000CD014095589EC0014D0A8E00CF09CE08AF009ED000005C950D015D004D0A" ;
	    attribute INIT_0A of bram : label is "00000000000000000000000000000000409EC003400A0080CF09CE08AF008E01" ;
	    attribute INIT_0B of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_0C of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_0D of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_0E of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_0F of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_10 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_11 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_12 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_13 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_14 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_15 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_16 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_17 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_18 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_19 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_1A of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_1B of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_1C of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_1D of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_1E of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_1F of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_20 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_21 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_22 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_23 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_24 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_25 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_26 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_27 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_28 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_29 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_2A of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_2B of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_2C of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_2D of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_2E of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_2F of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_30 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_31 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_32 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_33 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_34 of bram : label is "6961570E0A0D312E3076206E6F7275654E204C4448562048481667736D450502" ;
	    attribute INIT_35 of bram : label is "000000000000000000000000000000000000000000000A0D2E2E2E20676E6974" ;
	    attribute INIT_36 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_37 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_38 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_39 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_3A of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_3B of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_3C of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_3D of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_3E of bram : label is "4F13CF1303F81EF003F810100100000000000000000000000000000000000000" ;
	    attribute INIT_3F of bram : label is "8001A0004F10CF104F0353F82F014F0240005FEA51004109CF0B03F8CF0A9FE0" ;
	    attribute INITP_00 of bram : label is "E634A34E634ED2C8BFB4B22F4B22FEE22D2C8BED3D7FE9035FFA40FF3777777C" ;
	    attribute INITP_01 of bram : label is "00000000000000000000000000000000000000000000E3A59F4694C4683A33B4" ;
	    attribute INITP_02 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INITP_03 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INITP_04 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INITP_05 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INITP_06 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INITP_07 of bram : label is "E234F4B92CC00000000000000000000000000000000000000000000000000000" ;
	begin
	    bram : component RAMB16_S9_S18
	        generic map (
	            INIT_00 => X"000054024044501340545033405250464050505D404C5084404D0072008B0001",
	            INIT_01 => X"A1008001002F002F002F002FC2BAC0B99210028001000000006A40020080008B",
	            INIT_02 => X"0FFF40025C23E100C001002F002F002F002FC2BAC0B99210028001FF00FE5C16",
	            INIT_03 => X"4110C010007292004010C01000724213C2134210C01000720078A0005C30CF01",
	            INIT_04 => X"91004010C01000724113C1134110C010007200784002C27F006AC17E4113C113",
	            INIT_05 => X"C010007200784002D210006A92004010C01000724213C2134210C01000720078",
	            INIT_06 => X"400AC0034003506A200140024002C100006A91004010C01000724113C1134110",
	            INIT_07 => X"4078B0004F20CF034F0350782F014F02A000C0034003507220014002406AB000",
	            INIT_08 => X"8E00CE08CF090E800F0643E9C008C0090000008B0002006AA000548020024002",
	            INIT_09 => X"B000CD014095589EC0014D0A8E00CF09CE08AF009ED000005C950D015D004D0A",
	            INIT_0A => X"00000000000000000000000000000000409EC003400A0080CF09CE08AF008E01",
	            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_34 => X"6961570E0A0D312E3076206E6F7275654E204C4448562048481667736D450502",
	            INIT_35 => X"000000000000000000000000000000000000000000000A0D2E2E2E20676E6974",
	            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_3E => X"4F13CF1303F81EF003F810100100000000000000000000000000000000000000",
	            INIT_3F => X"8001A0004F10CF104F0353F82F014F0240005FEA51004109CF0B03F8CF0A9FE0",
	            INITP_00 => X"E634A34E634ED2C8BFB4B22F4B22FEE22D2C8BED3D7FE9035FFA40FF3777777C",
	            INITP_01 => X"00000000000000000000000000000000000000000000E3A59F4694C4683A33B4",
	            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INITP_07 => X"E234F4B92CC00000000000000000000000000000000000000000000000000000"
	        )
          
	        port map (
	            DIB   => "0000000000000000",
	            DIPB  => "00",
	            ENB   => '1',
	            WEB   => '0',
	            SSRB  => '0',
	            CLKB  => clk,
	            ADDRB => address,
	            DOB   => instruction( INSTSIZE - 3 downto 0 ),
	            DOPB  => instruction( INSTSIZE - 1 downto INSTSIZE - 2 ),
	            DIA   => ext_data( JDATASIZE - 2 downto 0 ),
	            DIPA  => ext_data( JDATASIZE - 1 downto JDATASIZE - 1 ),
	            ENA   => '1',
	            WEA   => ext_write,
	            SSRA  => '0',
	            CLKA  => clk,
	            ADDRA => ext_addr,
	            DOA   => out_data( JDATASIZE - 2 downto 0 ),
	            DOPA  => out_data( JDATASIZE - 1 downto JDATASIZE - 1 )
	        ) ;
	end generate ;

end architecture mix ;
