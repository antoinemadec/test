../../../multiple_cpu/src/noc.sv