../../../xorshift/src/cpu.sv