../../../multiple_cpu/src/cpu.sv